/*
  Eric Villasenor
  evillase@gmail.com

  interface to coordinate caches and
  implement coherence protocol
  TODO: make interface array of 2 and pass array, or something
*/
`ifndef CACHE_CONTROL_IF_VH
`define CACHE_CONTROL_IF_VH

// ram memory types
`include "cpu_types_pkg.vh"

// split this into cache_control_if and ram_if
interface cache_control_if;
  // import types
  import cpu_types_pkg::*;

  // access with cpuid on each processor
  parameter CPUS = 1;
  parameter CPUID = 0;

  // arbitration
  logic   [CPUS-1:0]       iwait, dwait, iREN, dREN, dWEN;
  word_t  [CPUS-1:0]       iload, dload, dstore;
  word_t  [CPUS-1:0]       iaddr, daddr;

  // coherence
  // CPUS = number of cpus parameter passed from system -> cc
  // ccwait         : lets a cache know it needs to block cpu
  // ccinv          : let a cache know it needs to invalidate entry
  // ccwrite        : high if cache is doing a write of addr
  // ccsnoopaddr    : the addr being sent to other cache with either (wb/inv)
  // cctrans        : high if the cache state is transitioning (i.e. I->S, I->M, etc...)
  logic   [CPUS-1:0]      ccwait, ccinv;
  logic   [CPUS-1:0]      ccwrite, cctrans;
  word_t  [CPUS-1:0]      ccsnoopaddr;

  // ram side
  logic                   ramWEN, ramREN;
  ramstate_t              ramstate;
  word_t                  ramaddr, ramstore, ramload;

  // controller ports to ram and caches
  modport cc (
            // cache inputs
    input   iREN, dREN, dWEN, dstore, iaddr, daddr,
            // ram inputs
            ramload, ramstate,
            // coherence inputs from cache
            ccwrite, cctrans,
            // cache outputs
    output  iwait, dwait, iload, dload,
            // ram outputs
            ramstore, ramaddr, ramWEN, ramREN,
            // coherence outputs to cache
            ccwait, ccinv, ccsnoopaddr
  );

  // icache ports to controller
  /*modport icache (
    input   iwait, iload,
    output  iREN, iaddr
  );

  // dcache ports to controller
  modport dcache (
    input   dwait, dload,
            ccwait, ccinv, ccsnoopaddr,
    output  dREN, dWEN, daddr, dstore,
            ccwrite, cctrans
<<<<<<< HEAD
=======
  );
  modport caches (
    input   iwait, iload, dwait, dload,
            ccwait, ccinv, ccsnoopaddr,
    output  iREN, iaddr, dREN, dWEN, daddr, dstore,
            ccwrite, cctrans
>>>>>>> 7dabfc3f11bbd03f1d249da3c2c0e8ce18ffaab5
  );
  modport caches (
    input   iwait, iload, dwait, dload,
            ccwait, ccinv, ccsnoopaddr,
    output  iREN, iaddr, dREN, dWEN, daddr, dstore,
            ccwrite, cctrans
  );*/

  modport caches (
    input   .iwait(iwait[CPUID]), 
    input   .iload(iload[CPUID]),
    input   .dwait(dwait[CPUID]), 
    input   .dload(dload[CPUID]),
    input   .ccwait(ccwait[CPUID]),
    input   .ccinv(ccinv[CPUID]),
    input   .ccsnoopaddr(ccsnoopaddr[CPUID]),

    output  .iREN(iREN[CPUID]),
    output  .iaddr(iaddr[CPUID]),
    output  .dREN(dREN[CPUID]),
    output  .dWEN(dWEN[CPUID]),
    output  .daddr(daddr[CPUID]),
    output  .dstore(dstore[CPUID]),
    output  .ccwrite(ccwrite[CPUID]),
    output  .cctrans(cctrans[CPUID])   
);

  modport icache (
    input   .iwait(iwait[CPUID]), 
    input   .iload(iload[CPUID]),

    output  .iREN(iREN[CPUID]),
    output  .iaddr(iaddr[CPUID])  
);

  modport icachetb (
    output   .iwait(iwait[CPUID]), 
    output   .iload(iload[CPUID]),

    input  .iREN(iREN[CPUID]),
    input  .iaddr(iaddr[CPUID])  
  );

  modport dcache (
    input   .dwait(dwait[CPUID]), 
    input   .dload(dload[CPUID]),
    input   .ccwait(ccwait[CPUID]),
    input   .ccinv(ccinv[CPUID]),
    input   .ccsnoopaddr(ccsnoopaddr[CPUID]),

    output  .dREN(dREN[CPUID]),
    output  .dWEN(dWEN[CPUID]),
    output  .daddr(daddr[CPUID]),
    output  .dstore(dstore[CPUID]),
    output  .ccwrite(ccwrite[CPUID]),
    output  .cctrans(cctrans[CPUID])   
);

  modport dcachetb (
    output   .dwait(dwait[CPUID]), 
    output   .dload(dload[CPUID]),
    output   .ccwait(ccwait[CPUID]),
    output   .ccinv(ccinv[CPUID]),
    output   .ccsnoopaddr(ccsnoopaddr[CPUID]),

    input  .dREN(dREN[CPUID]),
    input  .dWEN(dWEN[CPUID]),
    input  .daddr(daddr[CPUID]),
    input  .dstore(dstore[CPUID]),
    input  .ccwrite(ccwrite[CPUID]),
    input  .cctrans(cctrans[CPUID])   
  );



endinterface

`endif //CACHE_CONTROL_IF_VH
